
module CPU_Nios (
	clk_clk,
	leds_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	leds_export;
	input		reset_reset_n;
endmodule
