// CPU_Nios.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU_Nios (
		input  wire       clk_clk,       //   clk.clk
		output wire [7:0] leds_export,   //  leds.export
		input  wire       reset_reset_n  // reset.reset_n
	);

	wire  [31:0] cpu_nios_data_master_readdata;                          // mm_interconnect_0:cpu_Nios_data_master_readdata -> cpu_Nios:d_readdata
	wire         cpu_nios_data_master_waitrequest;                       // mm_interconnect_0:cpu_Nios_data_master_waitrequest -> cpu_Nios:d_waitrequest
	wire         cpu_nios_data_master_debugaccess;                       // cpu_Nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_Nios_data_master_debugaccess
	wire  [13:0] cpu_nios_data_master_address;                           // cpu_Nios:d_address -> mm_interconnect_0:cpu_Nios_data_master_address
	wire   [3:0] cpu_nios_data_master_byteenable;                        // cpu_Nios:d_byteenable -> mm_interconnect_0:cpu_Nios_data_master_byteenable
	wire         cpu_nios_data_master_read;                              // cpu_Nios:d_read -> mm_interconnect_0:cpu_Nios_data_master_read
	wire         cpu_nios_data_master_write;                             // cpu_Nios:d_write -> mm_interconnect_0:cpu_Nios_data_master_write
	wire  [31:0] cpu_nios_data_master_writedata;                         // cpu_Nios:d_writedata -> mm_interconnect_0:cpu_Nios_data_master_writedata
	wire  [31:0] cpu_nios_instruction_master_readdata;                   // mm_interconnect_0:cpu_Nios_instruction_master_readdata -> cpu_Nios:i_readdata
	wire         cpu_nios_instruction_master_waitrequest;                // mm_interconnect_0:cpu_Nios_instruction_master_waitrequest -> cpu_Nios:i_waitrequest
	wire  [13:0] cpu_nios_instruction_master_address;                    // cpu_Nios:i_address -> mm_interconnect_0:cpu_Nios_instruction_master_address
	wire         cpu_nios_instruction_master_read;                       // cpu_Nios:i_read -> mm_interconnect_0:cpu_Nios_instruction_master_read
	wire  [31:0] mm_interconnect_0_cpu_nios_debug_mem_slave_readdata;    // cpu_Nios:debug_mem_slave_readdata -> mm_interconnect_0:cpu_Nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_waitrequest; // cpu_Nios:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_Nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_debugaccess; // mm_interconnect_0:cpu_Nios_debug_mem_slave_debugaccess -> cpu_Nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_nios_debug_mem_slave_address;     // mm_interconnect_0:cpu_Nios_debug_mem_slave_address -> cpu_Nios:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_read;        // mm_interconnect_0:cpu_Nios_debug_mem_slave_read -> cpu_Nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_nios_debug_mem_slave_byteenable;  // mm_interconnect_0:cpu_Nios_debug_mem_slave_byteenable -> cpu_Nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_nios_debug_mem_slave_write;       // mm_interconnect_0:cpu_Nios_debug_mem_slave_write -> cpu_Nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_nios_debug_mem_slave_writedata;   // mm_interconnect_0:cpu_Nios_debug_mem_slave_writedata -> cpu_Nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_pio_s1_chipselect;                    // mm_interconnect_0:pio_s1_chipselect -> pio:chipselect
	wire  [31:0] mm_interconnect_0_pio_s1_readdata;                      // pio:readdata -> mm_interconnect_0:pio_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_s1_address;                       // mm_interconnect_0:pio_s1_address -> pio:address
	wire         mm_interconnect_0_pio_s1_write;                         // mm_interconnect_0:pio_s1_write -> pio:write_n
	wire  [31:0] mm_interconnect_0_pio_s1_writedata;                     // mm_interconnect_0:pio_s1_writedata -> pio:writedata
	wire         mm_interconnect_0_memory_ram_s1_chipselect;             // mm_interconnect_0:memory_RAM_s1_chipselect -> memory_RAM:chipselect
	wire  [31:0] mm_interconnect_0_memory_ram_s1_readdata;               // memory_RAM:readdata -> mm_interconnect_0:memory_RAM_s1_readdata
	wire   [9:0] mm_interconnect_0_memory_ram_s1_address;                // mm_interconnect_0:memory_RAM_s1_address -> memory_RAM:address
	wire   [3:0] mm_interconnect_0_memory_ram_s1_byteenable;             // mm_interconnect_0:memory_RAM_s1_byteenable -> memory_RAM:byteenable
	wire         mm_interconnect_0_memory_ram_s1_write;                  // mm_interconnect_0:memory_RAM_s1_write -> memory_RAM:write
	wire  [31:0] mm_interconnect_0_memory_ram_s1_writedata;              // mm_interconnect_0:memory_RAM_s1_writedata -> memory_RAM:writedata
	wire         mm_interconnect_0_memory_ram_s1_clken;                  // mm_interconnect_0:memory_RAM_s1_clken -> memory_RAM:clken
	wire         irq_mapper_receiver0_irq;                               // timer_interruption:irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_nios_irq_irq;                                       // irq_mapper:sender_irq -> cpu_Nios:irq
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [cpu_Nios:reset_n, irq_mapper:reset, memory_RAM:reset, mm_interconnect_0:cpu_Nios_reset_reset_bridge_in_reset_reset, pio:reset_n, rst_translator:in_reset, timer_interruption:reset_n]
	wire         rst_controller_reset_out_reset_req;                     // rst_controller:reset_req -> [cpu_Nios:reset_req, memory_RAM:reset_req, rst_translator:reset_req_in]

	CPU_Nios_cpu_Nios cpu_nios (
		.clk                                 (clk_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (cpu_nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_nios_data_master_read),                              //                          .read
		.d_readdata                          (cpu_nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_nios_data_master_write),                             //                          .write
		.d_writedata                         (cpu_nios_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_nios_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_nios_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                       //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	CPU_Nios_memory_RAM memory_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_memory_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	CPU_Nios_pio pio (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                          // external_connection.export
	);

	CPU_Nios_timer_interruption timer_interruption (
		.clk        (clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset), // reset.reset_n
		.address    (),                                //    s1.address
		.writedata  (),                                //      .writedata
		.readdata   (),                                //      .readdata
		.chipselect (),                                //      .chipselect
		.write_n    (),                                //      .write_n
		.irq        (irq_mapper_receiver0_irq)         //   irq.irq
	);

	CPU_Nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_cpu_clk_clk                            (clk_clk),                                                //                          clk_cpu_clk.clk
		.cpu_Nios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                         // cpu_Nios_reset_reset_bridge_in_reset.reset
		.cpu_Nios_data_master_address               (cpu_nios_data_master_address),                           //                 cpu_Nios_data_master.address
		.cpu_Nios_data_master_waitrequest           (cpu_nios_data_master_waitrequest),                       //                                     .waitrequest
		.cpu_Nios_data_master_byteenable            (cpu_nios_data_master_byteenable),                        //                                     .byteenable
		.cpu_Nios_data_master_read                  (cpu_nios_data_master_read),                              //                                     .read
		.cpu_Nios_data_master_readdata              (cpu_nios_data_master_readdata),                          //                                     .readdata
		.cpu_Nios_data_master_write                 (cpu_nios_data_master_write),                             //                                     .write
		.cpu_Nios_data_master_writedata             (cpu_nios_data_master_writedata),                         //                                     .writedata
		.cpu_Nios_data_master_debugaccess           (cpu_nios_data_master_debugaccess),                       //                                     .debugaccess
		.cpu_Nios_instruction_master_address        (cpu_nios_instruction_master_address),                    //          cpu_Nios_instruction_master.address
		.cpu_Nios_instruction_master_waitrequest    (cpu_nios_instruction_master_waitrequest),                //                                     .waitrequest
		.cpu_Nios_instruction_master_read           (cpu_nios_instruction_master_read),                       //                                     .read
		.cpu_Nios_instruction_master_readdata       (cpu_nios_instruction_master_readdata),                   //                                     .readdata
		.cpu_Nios_debug_mem_slave_address           (mm_interconnect_0_cpu_nios_debug_mem_slave_address),     //             cpu_Nios_debug_mem_slave.address
		.cpu_Nios_debug_mem_slave_write             (mm_interconnect_0_cpu_nios_debug_mem_slave_write),       //                                     .write
		.cpu_Nios_debug_mem_slave_read              (mm_interconnect_0_cpu_nios_debug_mem_slave_read),        //                                     .read
		.cpu_Nios_debug_mem_slave_readdata          (mm_interconnect_0_cpu_nios_debug_mem_slave_readdata),    //                                     .readdata
		.cpu_Nios_debug_mem_slave_writedata         (mm_interconnect_0_cpu_nios_debug_mem_slave_writedata),   //                                     .writedata
		.cpu_Nios_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_nios_debug_mem_slave_byteenable),  //                                     .byteenable
		.cpu_Nios_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_nios_debug_mem_slave_waitrequest), //                                     .waitrequest
		.cpu_Nios_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_nios_debug_mem_slave_debugaccess), //                                     .debugaccess
		.memory_RAM_s1_address                      (mm_interconnect_0_memory_ram_s1_address),                //                        memory_RAM_s1.address
		.memory_RAM_s1_write                        (mm_interconnect_0_memory_ram_s1_write),                  //                                     .write
		.memory_RAM_s1_readdata                     (mm_interconnect_0_memory_ram_s1_readdata),               //                                     .readdata
		.memory_RAM_s1_writedata                    (mm_interconnect_0_memory_ram_s1_writedata),              //                                     .writedata
		.memory_RAM_s1_byteenable                   (mm_interconnect_0_memory_ram_s1_byteenable),             //                                     .byteenable
		.memory_RAM_s1_chipselect                   (mm_interconnect_0_memory_ram_s1_chipselect),             //                                     .chipselect
		.memory_RAM_s1_clken                        (mm_interconnect_0_memory_ram_s1_clken),                  //                                     .clken
		.pio_s1_address                             (mm_interconnect_0_pio_s1_address),                       //                               pio_s1.address
		.pio_s1_write                               (mm_interconnect_0_pio_s1_write),                         //                                     .write
		.pio_s1_readdata                            (mm_interconnect_0_pio_s1_readdata),                      //                                     .readdata
		.pio_s1_writedata                           (mm_interconnect_0_pio_s1_writedata),                     //                                     .writedata
		.pio_s1_chipselect                          (mm_interconnect_0_pio_s1_chipselect)                     //                                     .chipselect
	);

	CPU_Nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_nios_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
