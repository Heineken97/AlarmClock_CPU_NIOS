// CPU_Nios_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU_Nios_tb (
	);

	wire        cpu_nios_inst_clk_bfm_clk_clk;       // CPU_Nios_inst_clk_bfm:clk -> [CPU_Nios_inst:clk_clk, CPU_Nios_inst_reset_bfm:clk]
	wire  [7:0] cpu_nios_inst_leds_export;           // CPU_Nios_inst:leds_export -> CPU_Nios_inst_leds_bfm:sig_export
	wire        cpu_nios_inst_reset_bfm_reset_reset; // CPU_Nios_inst_reset_bfm:reset -> CPU_Nios_inst:reset_reset_n

	CPU_Nios cpu_nios_inst (
		.clk_clk       (cpu_nios_inst_clk_bfm_clk_clk),       //   clk.clk
		.leds_export   (cpu_nios_inst_leds_export),           //  leds.export
		.reset_reset_n (cpu_nios_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) cpu_nios_inst_clk_bfm (
		.clk (cpu_nios_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm cpu_nios_inst_leds_bfm (
		.sig_export (cpu_nios_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) cpu_nios_inst_reset_bfm (
		.reset (cpu_nios_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (cpu_nios_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
